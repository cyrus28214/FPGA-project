`timescale 1ns/1ps

module music_player(
    input clk, // 100 MHz
    output beep
);

reg [31:0] i, p, cnt;
parameter MAXN = 150;
reg [31:0] pos[MAXN-1:0];
reg [7:0] note[MAXN-1:0];
initial begin
    note[0] = 76;
    note[1] = 71;
    note[2] = 69;
    note[3] = 72;
    note[4] = 68;
    note[5] = 0;
    note[6] = 71;
    note[7] = 69;
    note[8] = 57;
    note[9] = 64;
    note[10] = 65;
    note[11] = 0;
    note[12] = 76;
    note[13] = 71;
    note[14] = 69;
    note[15] = 72;
    note[16] = 68;
    note[17] = 0;
    note[18] = 71;
    note[19] = 69;
    note[20] = 57;
    note[21] = 64;
    note[22] = 65;
    note[23] = 0;
    note[24] = 76;
    note[25] = 69;
    note[26] = 65;
    note[27] = 67;
    note[28] = 62;
    note[29] = 64;
    note[30] = 0;
    note[31] = 76;
    note[32] = 69;
    note[33] = 65;
    note[34] = 67;
    note[35] = 74;
    note[36] = 72;
    note[37] = 70;
    note[38] = 69;
    note[39] = 0;
    note[40] = 69;
    note[41] = 71;
    note[42] = 72;
    note[43] = 0;
    note[44] = 72;
    note[45] = 74;
    note[46] = 76;
    note[47] = 0;
    note[48] = 71;
    note[49] = 64;
    note[50] = 0;
    note[51] = 76;
    note[52] = 0;
    note[53] = 62;
    note[54] = 0;
    note[55] = 62;
    note[56] = 64;
    note[57] = 69;
    note[58] = 62;
    note[59] = 64;
    note[60] = 69;
    note[61] = 70;
    note[62] = 62;
    note[63] = 64;
    note[64] = 70;
    note[65] = 69;
    note[66] = 0;
    note[67] = 62;
    note[68] = 64;
    note[69] = 69;
    note[70] = 62;
    note[71] = 64;
    note[72] = 69;
    note[73] = 67;
    note[74] = 62;
    note[75] = 64;
    note[76] = 67;
    note[77] = 69;
    note[78] = 0;
    note[79] = 62;
    note[80] = 64;
    note[81] = 69;
    note[82] = 62;
    note[83] = 64;
    note[84] = 69;
    note[85] = 70;
    note[86] = 62;
    note[87] = 64;
    note[88] = 70;
    note[89] = 69;
    note[90] = 0;
    note[91] = 62;
    note[92] = 64;
    note[93] = 69;
    note[94] = 62;
    note[95] = 64;
    note[96] = 69;
    note[97] = 67;
    note[98] = 62;
    note[99] = 64;
    note[100] = 67;
    note[101] = 76;
    note[102] = 74;
    note[103] = 69;
    note[104] = 71;
    note[105] = 62;
    note[106] = 69;
    note[107] = 71;
    note[108] = 74;
    note[109] = 76;
    note[110] = 74;
    note[111] = 76;
    note[112] = 0;
    note[113] = 76;
    note[114] = 0;
    note[115] = 76;
    note[116] = 74;
    note[117] = 69;
    note[118] = 71;
    note[119] = 62;
    note[120] = 69;
    note[121] = 71;
    note[122] = 74;
    note[123] = 76;
    note[124] = 71;
    note[125] = 74;
    note[126] = 76;
    note[127] = 0;
    note[128] = 76;
    note[129] = 81;
    note[130] = 83;
    note[131] = 76;
    note[132] = 0;
    note[133] = 64;
    note[134] = 0;
    note[135] = 72;
    note[136] = 74;
    note[137] = 76;
    note[138] = 83;
    note[139] = 81;
    note[140] = 76;
    note[141] = 74;
    note[142] = 76;
    note[143] = 69;
    note[144] = 71;
    note[145] = 72;
    note[146] = 74;
    note[147] = 71;
    note[148] = 0;
    note[149] = 76;
end
initial begin
    pos[0] = 500;
    pos[1] = 1000;
    pos[2] = 1500;
    pos[3] = 2000;
    pos[4] = 2500;
    pos[5] = 3000;
    pos[6] = 3500;
    pos[7] = 4000;
    pos[8] = 4500;
    pos[9] = 5000;
    pos[10] = 5500;
    pos[11] = 6000;
    pos[12] = 6500;
    pos[13] = 7000;
    pos[14] = 7500;
    pos[15] = 8000;
    pos[16] = 8500;
    pos[17] = 9000;
    pos[18] = 9500;
    pos[19] = 10000;
    pos[20] = 10500;
    pos[21] = 11000;
    pos[22] = 11500;
    pos[23] = 12000;
    pos[24] = 12500;
    pos[25] = 13000;
    pos[26] = 13500;
    pos[27] = 14500;
    pos[28] = 15000;
    pos[29] = 17750;
    pos[30] = 18125;
    pos[31] = 18625;
    pos[32] = 19125;
    pos[33] = 19625;
    pos[34] = 20625;
    pos[35] = 21125;
    pos[36] = 23125;
    pos[37] = 24125;
    pos[38] = 25875;
    pos[39] = 26125;
    pos[40] = 26625;
    pos[41] = 27125;
    pos[42] = 29000;
    pos[43] = 29125;
    pos[44] = 29625;
    pos[45] = 30125;
    pos[46] = 32000;
    pos[47] = 32250;
    pos[48] = 33250;
    pos[49] = 36000;
    pos[50] = 36250;
    pos[51] = 36500;
    pos[52] = 36750;
    pos[53] = 37000;
    pos[54] = 36750;
    pos[55] = 37000;
    pos[56] = 37250;
    pos[57] = 37500;
    pos[58] = 37750;
    pos[59] = 38000;
    pos[60] = 38250;
    pos[61] = 38500;
    pos[62] = 38750;
    pos[63] = 39000;
    pos[64] = 39250;
    pos[65] = 39625;
    pos[66] = 39750;
    pos[67] = 40000;
    pos[68] = 40250;
    pos[69] = 40500;
    pos[70] = 40750;
    pos[71] = 41000;
    pos[72] = 41250;
    pos[73] = 41500;
    pos[74] = 41750;
    pos[75] = 42000;
    pos[76] = 42250;
    pos[77] = 42500;
    pos[78] = 42750;
    pos[79] = 43000;
    pos[80] = 43250;
    pos[81] = 43500;
    pos[82] = 43750;
    pos[83] = 44000;
    pos[84] = 44250;
    pos[85] = 44500;
    pos[86] = 44750;
    pos[87] = 45000;
    pos[88] = 45250;
    pos[89] = 45500;
    pos[90] = 45750;
    pos[91] = 46000;
    pos[92] = 46250;
    pos[93] = 46500;
    pos[94] = 46750;
    pos[95] = 47000;
    pos[96] = 47250;
    pos[97] = 47500;
    pos[98] = 47750;
    pos[99] = 48000;
    pos[100] = 48250;
    pos[101] = 48500;
    pos[102] = 48750;
    pos[103] = 49000;
    pos[104] = 49250;
    pos[105] = 49500;
    pos[106] = 49750;
    pos[107] = 50000;
    pos[108] = 50250;
    pos[109] = 50500;
    pos[110] = 50750;
    pos[111] = 50947;
    pos[112] = 51000;
    pos[113] = 51083;
    pos[114] = 51250;
    pos[115] = 51500;
    pos[116] = 51750;
    pos[117] = 52000;
    pos[118] = 52250;
    pos[119] = 52500;
    pos[120] = 52750;
    pos[121] = 53000;
    pos[122] = 53250;
    pos[123] = 53500;
    pos[124] = 53750;
    pos[125] = 54000;
    pos[126] = 54234;
    pos[127] = 54250;
    pos[128] = 55250;
    pos[129] = 56250;
    pos[130] = 57250;
    pos[131] = 58625;
    pos[132] = 59250;
    pos[133] = 60250;
    pos[134] = 60375;
    pos[135] = 60875;
    pos[136] = 61375;
    pos[137] = 61875;
    pos[138] = 62375;
    pos[139] = 62875;
    pos[140] = 63375;
    pos[141] = 63875;
    pos[142] = 64375;
    pos[143] = 64875;
    pos[144] = 65375;
    pos[145] = 65875;
    pos[146] = 66375;
    pos[147] = 71875;
    pos[148] = 75875;
    pos[149] = 75901;
end


wire clk_out;
clk_1ms getClk(
    .clk(clk),
    .clk_1ms(clk_out)
);

initial begin
    cnt = 0;
    p = 0;
end

always @(posedge clk_out) begin
    if( cnt >= pos[MAXN-1] ) begin
        cnt <= 0;
        p <= 0;
    end else begin
        cnt <= cnt + 1;
        p <= pos[p] <= cnt ? p + 1 : p;
    end
end

wire [7:0] note_in = note[p];
buzzer inst(
    .clk(clk),
    .note(note_in),
    .beep(beep)
);

endmodule